module src;
endmodule: src